module MIPS_single_cycle #(parameter depth = 1024, width = 8)(
    input           wire                                   clk,
    input           wire                                   rst,
    input           wire      [$clog2(depth)-1:0]          instr_MEM_write_address,
    input           wire                                   instr_MEM_WE,
    
    

);
    
endmodule