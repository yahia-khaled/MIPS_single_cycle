module INST_MEM #(parameter depth = 1100, width = 8) (
    input       wire            [4*width-1:0]             Read_address,
    output      wire            [4*width-1:0]              RD
);


(* rom_style = "block" *)  // Force Vivado to infer Block RAM (BRAM)
reg     [width-1:0]       MEM     [0:depth-1];

assign RD = {MEM[Read_address+3], MEM[Read_address+2], MEM[Read_address+1], MEM[Read_address]};


integer i;

initial begin
    MEM[0] = 8'hfc;
    MEM[1] = 8'h7f;
    MEM[2] = 8'h1d;
    MEM[3] = 8'h20;
    MEM[4] = 8'h80;
    MEM[5] = 8'h10;
    MEM[6] = 8'h1c;
    MEM[7] = 8'h20;
    MEM[8] = 8'h00;
    MEM[9] = 8'h01;
    MEM[10] = 8'h00;
    MEM[11] = 8'h0c;
    MEM[12] = 8'h00;
    MEM[13] = 8'h00;
    MEM[14] = 8'h00;
    MEM[15] = 8'h00;
    MEM[16] = 8'h00;
    MEM[17] = 8'h00;
    MEM[18] = 8'h00;
    MEM[19] = 8'h00;
    MEM[20] = 8'h00;
    MEM[21] = 8'h00;
    MEM[22] = 8'h00;
    MEM[23] = 8'h00;
    MEM[24] = 8'h00;
    MEM[25] = 8'h00;
    MEM[26] = 8'h00;
    MEM[27] = 8'h00;
    MEM[28] = 8'h00;
    MEM[29] = 8'h00;
    MEM[30] = 8'h00;
    MEM[31] = 8'h00;
    MEM[32] = 8'h00;
    MEM[33] = 8'h00;
    MEM[34] = 8'h00;
    MEM[35] = 8'h00;
    MEM[36] = 8'h00;
    MEM[37] = 8'h00;
    MEM[38] = 8'h00;
    MEM[39] = 8'h00;
    MEM[40] = 8'h00;
    MEM[41] = 8'h00;
    MEM[42] = 8'h00;
    MEM[43] = 8'h00;
    MEM[44] = 8'h00;
    MEM[45] = 8'h00;
    MEM[46] = 8'h00;
    MEM[47] = 8'h00;
    MEM[48] = 8'h00;
    MEM[49] = 8'h00;
    MEM[50] = 8'h00;
    MEM[51] = 8'h00;
    MEM[52] = 8'h00;
    MEM[53] = 8'h00;
    MEM[54] = 8'h00;
    MEM[55] = 8'h00;
    MEM[56] = 8'h00;
    MEM[57] = 8'h00;
    MEM[58] = 8'h00;
    MEM[59] = 8'h00;
    MEM[60] = 8'h00;
    MEM[61] = 8'h00;
    MEM[62] = 8'h00;
    MEM[63] = 8'h00;
    MEM[64] = 8'h00;
    MEM[65] = 8'h00;
    MEM[66] = 8'h00;
    MEM[67] = 8'h00;
    MEM[68] = 8'h00;
    MEM[69] = 8'h00;
    MEM[70] = 8'h00;
    MEM[71] = 8'h00;
    MEM[72] = 8'h00;
    MEM[73] = 8'h00;
    MEM[74] = 8'h00;
    MEM[75] = 8'h00;
    MEM[76] = 8'h00;
    MEM[77] = 8'h00;
    MEM[78] = 8'h00;
    MEM[79] = 8'h00;
    MEM[80] = 8'h00;
    MEM[81] = 8'h00;
    MEM[82] = 8'h00;
    MEM[83] = 8'h00;
    MEM[84] = 8'h00;
    MEM[85] = 8'h00;
    MEM[86] = 8'h00;
    MEM[87] = 8'h00;
    MEM[88] = 8'h00;
    MEM[89] = 8'h00;
    MEM[90] = 8'h00;
    MEM[91] = 8'h00;
    MEM[92] = 8'h00;
    MEM[93] = 8'h00;
    MEM[94] = 8'h00;
    MEM[95] = 8'h00;
    MEM[96] = 8'h00;
    MEM[97] = 8'h00;
    MEM[98] = 8'h00;
    MEM[99] = 8'h00;
    MEM[100] = 8'h00;
    MEM[101] = 8'h00;
    MEM[102] = 8'h00;
    MEM[103] = 8'h00;
    MEM[104] = 8'h00;
    MEM[105] = 8'h00;
    MEM[106] = 8'h00;
    MEM[107] = 8'h00;
    MEM[108] = 8'h00;
    MEM[109] = 8'h00;
    MEM[110] = 8'h00;
    MEM[111] = 8'h00;
    MEM[112] = 8'h00;
    MEM[113] = 8'h00;
    MEM[114] = 8'h00;
    MEM[115] = 8'h00;
    MEM[116] = 8'h00;
    MEM[117] = 8'h00;
    MEM[118] = 8'h00;
    MEM[119] = 8'h00;
    MEM[120] = 8'h00;
    MEM[121] = 8'h00;
    MEM[122] = 8'h00;
    MEM[123] = 8'h00;
    MEM[124] = 8'h00;
    MEM[125] = 8'h00;
    MEM[126] = 8'h00;
    MEM[127] = 8'h00;
    MEM[128] = 8'h00;
    MEM[129] = 8'h00;
    MEM[130] = 8'h00;
    MEM[131] = 8'h00;
    MEM[132] = 8'h00;
    MEM[133] = 8'h00;
    MEM[134] = 8'h00;
    MEM[135] = 8'h00;
    MEM[136] = 8'h00;
    MEM[137] = 8'h00;
    MEM[138] = 8'h00;
    MEM[139] = 8'h00;
    MEM[140] = 8'h00;
    MEM[141] = 8'h00;
    MEM[142] = 8'h00;
    MEM[143] = 8'h00;
    MEM[144] = 8'h00;
    MEM[145] = 8'h00;
    MEM[146] = 8'h00;
    MEM[147] = 8'h00;
    MEM[148] = 8'h00;
    MEM[149] = 8'h00;
    MEM[150] = 8'h00;
    MEM[151] = 8'h00;
    MEM[152] = 8'h00;
    MEM[153] = 8'h00;
    MEM[154] = 8'h00;
    MEM[155] = 8'h00;
    MEM[156] = 8'h00;
    MEM[157] = 8'h00;
    MEM[158] = 8'h00;
    MEM[159] = 8'h00;
    MEM[160] = 8'h00;
    MEM[161] = 8'h00;
    MEM[162] = 8'h00;
    MEM[163] = 8'h00;
    MEM[164] = 8'h00;
    MEM[165] = 8'h00;
    MEM[166] = 8'h00;
    MEM[167] = 8'h00;
    MEM[168] = 8'h00;
    MEM[169] = 8'h00;
    MEM[170] = 8'h00;
    MEM[171] = 8'h00;
    MEM[172] = 8'h00;
    MEM[173] = 8'h00;
    MEM[174] = 8'h00;
    MEM[175] = 8'h00;
    MEM[176] = 8'h00;
    MEM[177] = 8'h00;
    MEM[178] = 8'h00;
    MEM[179] = 8'h00;
    MEM[180] = 8'h00;
    MEM[181] = 8'h00;
    MEM[182] = 8'h00;
    MEM[183] = 8'h00;
    MEM[184] = 8'h00;
    MEM[185] = 8'h00;
    MEM[186] = 8'h00;
    MEM[187] = 8'h00;
    MEM[188] = 8'h00;
    MEM[189] = 8'h00;
    MEM[190] = 8'h00;
    MEM[191] = 8'h00;
    MEM[192] = 8'h00;
    MEM[193] = 8'h00;
    MEM[194] = 8'h00;
    MEM[195] = 8'h00;
    MEM[196] = 8'h00;
    MEM[197] = 8'h00;
    MEM[198] = 8'h00;
    MEM[199] = 8'h00;
    MEM[200] = 8'h00;
    MEM[201] = 8'h00;
    MEM[202] = 8'h00;
    MEM[203] = 8'h00;
    MEM[204] = 8'h00;
    MEM[205] = 8'h00;
    MEM[206] = 8'h00;
    MEM[207] = 8'h00;
    MEM[208] = 8'h00;
    MEM[209] = 8'h00;
    MEM[210] = 8'h00;
    MEM[211] = 8'h00;
    MEM[212] = 8'h00;
    MEM[213] = 8'h00;
    MEM[214] = 8'h00;
    MEM[215] = 8'h00;
    MEM[216] = 8'h00;
    MEM[217] = 8'h00;
    MEM[218] = 8'h00;
    MEM[219] = 8'h00;
    MEM[220] = 8'h00;
    MEM[221] = 8'h00;
    MEM[222] = 8'h00;
    MEM[223] = 8'h00;
    MEM[224] = 8'h00;
    MEM[225] = 8'h00;
    MEM[226] = 8'h00;
    MEM[227] = 8'h00;
    MEM[228] = 8'h00;
    MEM[229] = 8'h00;
    MEM[230] = 8'h00;
    MEM[231] = 8'h00;
    MEM[232] = 8'h00;
    MEM[233] = 8'h00;
    MEM[234] = 8'h00;
    MEM[235] = 8'h00;
    MEM[236] = 8'h00;
    MEM[237] = 8'h00;
    MEM[238] = 8'h00;
    MEM[239] = 8'h00;
    MEM[240] = 8'h00;
    MEM[241] = 8'h00;
    MEM[242] = 8'h00;
    MEM[243] = 8'h00;
    MEM[244] = 8'h00;
    MEM[245] = 8'h00;
    MEM[246] = 8'h00;
    MEM[247] = 8'h00;
    MEM[248] = 8'h00;
    MEM[249] = 8'h00;
    MEM[250] = 8'h00;
    MEM[251] = 8'h00;
    MEM[252] = 8'h00;
    MEM[253] = 8'h00;
    MEM[254] = 8'h00;
    MEM[255] = 8'h00;
    MEM[256] = 8'h00;
    MEM[257] = 8'h00;
    MEM[258] = 8'h00;
    MEM[259] = 8'h00;
    MEM[260] = 8'h00;
    MEM[261] = 8'h00;
    MEM[262] = 8'h00;
    MEM[263] = 8'h00;
    MEM[264] = 8'h00;
    MEM[265] = 8'h00;
    MEM[266] = 8'h00;
    MEM[267] = 8'h00;
    MEM[268] = 8'h00;
    MEM[269] = 8'h00;
    MEM[270] = 8'h00;
    MEM[271] = 8'h00;
    MEM[272] = 8'h00;
    MEM[273] = 8'h00;
    MEM[274] = 8'h00;
    MEM[275] = 8'h00;
    MEM[276] = 8'h00;
    MEM[277] = 8'h00;
    MEM[278] = 8'h00;
    MEM[279] = 8'h00;
    MEM[280] = 8'h00;
    MEM[281] = 8'h00;
    MEM[282] = 8'h00;
    MEM[283] = 8'h00;
    MEM[284] = 8'h00;
    MEM[285] = 8'h00;
    MEM[286] = 8'h00;
    MEM[287] = 8'h00;
    MEM[288] = 8'h00;
    MEM[289] = 8'h00;
    MEM[290] = 8'h00;
    MEM[291] = 8'h00;
    MEM[292] = 8'h00;
    MEM[293] = 8'h00;
    MEM[294] = 8'h00;
    MEM[295] = 8'h00;
    MEM[296] = 8'h00;
    MEM[297] = 8'h00;
    MEM[298] = 8'h00;
    MEM[299] = 8'h00;
    MEM[300] = 8'h00;
    MEM[301] = 8'h00;
    MEM[302] = 8'h00;
    MEM[303] = 8'h00;
    MEM[304] = 8'h00;
    MEM[305] = 8'h00;
    MEM[306] = 8'h00;
    MEM[307] = 8'h00;
    MEM[308] = 8'h00;
    MEM[309] = 8'h00;
    MEM[310] = 8'h00;
    MEM[311] = 8'h00;
    MEM[312] = 8'h00;
    MEM[313] = 8'h00;
    MEM[314] = 8'h00;
    MEM[315] = 8'h00;
    MEM[316] = 8'h00;
    MEM[317] = 8'h00;
    MEM[318] = 8'h00;
    MEM[319] = 8'h00;
    MEM[320] = 8'h00;
    MEM[321] = 8'h00;
    MEM[322] = 8'h00;
    MEM[323] = 8'h00;
    MEM[324] = 8'h00;
    MEM[325] = 8'h00;
    MEM[326] = 8'h00;
    MEM[327] = 8'h00;
    MEM[328] = 8'h00;
    MEM[329] = 8'h00;
    MEM[330] = 8'h00;
    MEM[331] = 8'h00;
    MEM[332] = 8'h00;
    MEM[333] = 8'h00;
    MEM[334] = 8'h00;
    MEM[335] = 8'h00;
    MEM[336] = 8'h00;
    MEM[337] = 8'h00;
    MEM[338] = 8'h00;
    MEM[339] = 8'h00;
    MEM[340] = 8'h00;
    MEM[341] = 8'h00;
    MEM[342] = 8'h00;
    MEM[343] = 8'h00;
    MEM[344] = 8'h00;
    MEM[345] = 8'h00;
    MEM[346] = 8'h00;
    MEM[347] = 8'h00;
    MEM[348] = 8'h00;
    MEM[349] = 8'h00;
    MEM[350] = 8'h00;
    MEM[351] = 8'h00;
    MEM[352] = 8'h00;
    MEM[353] = 8'h00;
    MEM[354] = 8'h00;
    MEM[355] = 8'h00;
    MEM[356] = 8'h00;
    MEM[357] = 8'h00;
    MEM[358] = 8'h00;
    MEM[359] = 8'h00;
    MEM[360] = 8'h00;
    MEM[361] = 8'h00;
    MEM[362] = 8'h00;
    MEM[363] = 8'h00;
    MEM[364] = 8'h00;
    MEM[365] = 8'h00;
    MEM[366] = 8'h00;
    MEM[367] = 8'h00;
    MEM[368] = 8'h00;
    MEM[369] = 8'h00;
    MEM[370] = 8'h00;
    MEM[371] = 8'h00;
    MEM[372] = 8'h00;
    MEM[373] = 8'h00;
    MEM[374] = 8'h00;
    MEM[375] = 8'h00;
    MEM[376] = 8'h00;
    MEM[377] = 8'h00;
    MEM[378] = 8'h00;
    MEM[379] = 8'h00;
    MEM[380] = 8'h00;
    MEM[381] = 8'h00;
    MEM[382] = 8'h00;
    MEM[383] = 8'h00;
    MEM[384] = 8'h00;
    MEM[385] = 8'h00;
    MEM[386] = 8'h00;
    MEM[387] = 8'h00;
    MEM[388] = 8'h00;
    MEM[389] = 8'h00;
    MEM[390] = 8'h00;
    MEM[391] = 8'h00;
    MEM[392] = 8'h00;
    MEM[393] = 8'h00;
    MEM[394] = 8'h00;
    MEM[395] = 8'h00;
    MEM[396] = 8'h00;
    MEM[397] = 8'h00;
    MEM[398] = 8'h00;
    MEM[399] = 8'h00;
    MEM[400] = 8'h00;
    MEM[401] = 8'h00;
    MEM[402] = 8'h00;
    MEM[403] = 8'h00;
    MEM[404] = 8'h00;
    MEM[405] = 8'h00;
    MEM[406] = 8'h00;
    MEM[407] = 8'h00;
    MEM[408] = 8'h00;
    MEM[409] = 8'h00;
    MEM[410] = 8'h00;
    MEM[411] = 8'h00;
    MEM[412] = 8'h00;
    MEM[413] = 8'h00;
    MEM[414] = 8'h00;
    MEM[415] = 8'h00;
    MEM[416] = 8'h00;
    MEM[417] = 8'h00;
    MEM[418] = 8'h00;
    MEM[419] = 8'h00;
    MEM[420] = 8'h00;
    MEM[421] = 8'h00;
    MEM[422] = 8'h00;
    MEM[423] = 8'h00;
    MEM[424] = 8'h00;
    MEM[425] = 8'h00;
    MEM[426] = 8'h00;
    MEM[427] = 8'h00;
    MEM[428] = 8'h00;
    MEM[429] = 8'h00;
    MEM[430] = 8'h00;
    MEM[431] = 8'h00;
    MEM[432] = 8'h00;
    MEM[433] = 8'h00;
    MEM[434] = 8'h00;
    MEM[435] = 8'h00;
    MEM[436] = 8'h00;
    MEM[437] = 8'h00;
    MEM[438] = 8'h00;
    MEM[439] = 8'h00;
    MEM[440] = 8'h00;
    MEM[441] = 8'h00;
    MEM[442] = 8'h00;
    MEM[443] = 8'h00;
    MEM[444] = 8'h00;
    MEM[445] = 8'h00;
    MEM[446] = 8'h00;
    MEM[447] = 8'h00;
    MEM[448] = 8'h00;
    MEM[449] = 8'h00;
    MEM[450] = 8'h00;
    MEM[451] = 8'h00;
    MEM[452] = 8'h00;
    MEM[453] = 8'h00;
    MEM[454] = 8'h00;
    MEM[455] = 8'h00;
    MEM[456] = 8'h00;
    MEM[457] = 8'h00;
    MEM[458] = 8'h00;
    MEM[459] = 8'h00;
    MEM[460] = 8'h00;
    MEM[461] = 8'h00;
    MEM[462] = 8'h00;
    MEM[463] = 8'h00;
    MEM[464] = 8'h00;
    MEM[465] = 8'h00;
    MEM[466] = 8'h00;
    MEM[467] = 8'h00;
    MEM[468] = 8'h00;
    MEM[469] = 8'h00;
    MEM[470] = 8'h00;
    MEM[471] = 8'h00;
    MEM[472] = 8'h00;
    MEM[473] = 8'h00;
    MEM[474] = 8'h00;
    MEM[475] = 8'h00;
    MEM[476] = 8'h00;
    MEM[477] = 8'h00;
    MEM[478] = 8'h00;
    MEM[479] = 8'h00;
    MEM[480] = 8'h00;
    MEM[481] = 8'h00;
    MEM[482] = 8'h00;
    MEM[483] = 8'h00;
    MEM[484] = 8'h00;
    MEM[485] = 8'h00;
    MEM[486] = 8'h00;
    MEM[487] = 8'h00;
    MEM[488] = 8'h00;
    MEM[489] = 8'h00;
    MEM[490] = 8'h00;
    MEM[491] = 8'h00;
    MEM[492] = 8'h00;
    MEM[493] = 8'h00;
    MEM[494] = 8'h00;
    MEM[495] = 8'h00;
    MEM[496] = 8'h00;
    MEM[497] = 8'h00;
    MEM[498] = 8'h00;
    MEM[499] = 8'h00;
    MEM[500] = 8'h00;
    MEM[501] = 8'h00;
    MEM[502] = 8'h00;
    MEM[503] = 8'h00;
    MEM[504] = 8'h00;
    MEM[505] = 8'h00;
    MEM[506] = 8'h00;
    MEM[507] = 8'h00;
    MEM[508] = 8'h00;
    MEM[509] = 8'h00;
    MEM[510] = 8'h00;
    MEM[511] = 8'h00;
    MEM[512] = 8'h00;
    MEM[513] = 8'h00;
    MEM[514] = 8'h00;
    MEM[515] = 8'h00;
    MEM[516] = 8'h00;
    MEM[517] = 8'h00;
    MEM[518] = 8'h00;
    MEM[519] = 8'h00;
    MEM[520] = 8'h00;
    MEM[521] = 8'h00;
    MEM[522] = 8'h00;
    MEM[523] = 8'h00;
    MEM[524] = 8'h00;
    MEM[525] = 8'h00;
    MEM[526] = 8'h00;
    MEM[527] = 8'h00;
    MEM[528] = 8'h00;
    MEM[529] = 8'h00;
    MEM[530] = 8'h00;
    MEM[531] = 8'h00;
    MEM[532] = 8'h00;
    MEM[533] = 8'h00;
    MEM[534] = 8'h00;
    MEM[535] = 8'h00;
    MEM[536] = 8'h00;
    MEM[537] = 8'h00;
    MEM[538] = 8'h00;
    MEM[539] = 8'h00;
    MEM[540] = 8'h00;
    MEM[541] = 8'h00;
    MEM[542] = 8'h00;
    MEM[543] = 8'h00;
    MEM[544] = 8'h00;
    MEM[545] = 8'h00;
    MEM[546] = 8'h00;
    MEM[547] = 8'h00;
    MEM[548] = 8'h00;
    MEM[549] = 8'h00;
    MEM[550] = 8'h00;
    MEM[551] = 8'h00;
    MEM[552] = 8'h00;
    MEM[553] = 8'h00;
    MEM[554] = 8'h00;
    MEM[555] = 8'h00;
    MEM[556] = 8'h00;
    MEM[557] = 8'h00;
    MEM[558] = 8'h00;
    MEM[559] = 8'h00;
    MEM[560] = 8'h00;
    MEM[561] = 8'h00;
    MEM[562] = 8'h00;
    MEM[563] = 8'h00;
    MEM[564] = 8'h00;
    MEM[565] = 8'h00;
    MEM[566] = 8'h00;
    MEM[567] = 8'h00;
    MEM[568] = 8'h00;
    MEM[569] = 8'h00;
    MEM[570] = 8'h00;
    MEM[571] = 8'h00;
    MEM[572] = 8'h00;
    MEM[573] = 8'h00;
    MEM[574] = 8'h00;
    MEM[575] = 8'h00;
    MEM[576] = 8'h00;
    MEM[577] = 8'h00;
    MEM[578] = 8'h00;
    MEM[579] = 8'h00;
    MEM[580] = 8'h00;
    MEM[581] = 8'h00;
    MEM[582] = 8'h00;
    MEM[583] = 8'h00;
    MEM[584] = 8'h00;
    MEM[585] = 8'h00;
    MEM[586] = 8'h00;
    MEM[587] = 8'h00;
    MEM[588] = 8'h00;
    MEM[589] = 8'h00;
    MEM[590] = 8'h00;
    MEM[591] = 8'h00;
    MEM[592] = 8'h00;
    MEM[593] = 8'h00;
    MEM[594] = 8'h00;
    MEM[595] = 8'h00;
    MEM[596] = 8'h00;
    MEM[597] = 8'h00;
    MEM[598] = 8'h00;
    MEM[599] = 8'h00;
    MEM[600] = 8'h00;
    MEM[601] = 8'h00;
    MEM[602] = 8'h00;
    MEM[603] = 8'h00;
    MEM[604] = 8'h00;
    MEM[605] = 8'h00;
    MEM[606] = 8'h00;
    MEM[607] = 8'h00;
    MEM[608] = 8'h00;
    MEM[609] = 8'h00;
    MEM[610] = 8'h00;
    MEM[611] = 8'h00;
    MEM[612] = 8'h00;
    MEM[613] = 8'h00;
    MEM[614] = 8'h00;
    MEM[615] = 8'h00;
    MEM[616] = 8'h00;
    MEM[617] = 8'h00;
    MEM[618] = 8'h00;
    MEM[619] = 8'h00;
    MEM[620] = 8'h00;
    MEM[621] = 8'h00;
    MEM[622] = 8'h00;
    MEM[623] = 8'h00;
    MEM[624] = 8'h00;
    MEM[625] = 8'h00;
    MEM[626] = 8'h00;
    MEM[627] = 8'h00;
    MEM[628] = 8'h00;
    MEM[629] = 8'h00;
    MEM[630] = 8'h00;
    MEM[631] = 8'h00;
    MEM[632] = 8'h00;
    MEM[633] = 8'h00;
    MEM[634] = 8'h00;
    MEM[635] = 8'h00;
    MEM[636] = 8'h00;
    MEM[637] = 8'h00;
    MEM[638] = 8'h00;
    MEM[639] = 8'h00;
    MEM[640] = 8'h00;
    MEM[641] = 8'h00;
    MEM[642] = 8'h00;
    MEM[643] = 8'h00;
    MEM[644] = 8'h00;
    MEM[645] = 8'h00;
    MEM[646] = 8'h00;
    MEM[647] = 8'h00;
    MEM[648] = 8'h00;
    MEM[649] = 8'h00;
    MEM[650] = 8'h00;
    MEM[651] = 8'h00;
    MEM[652] = 8'h00;
    MEM[653] = 8'h00;
    MEM[654] = 8'h00;
    MEM[655] = 8'h00;
    MEM[656] = 8'h00;
    MEM[657] = 8'h00;
    MEM[658] = 8'h00;
    MEM[659] = 8'h00;
    MEM[660] = 8'h00;
    MEM[661] = 8'h00;
    MEM[662] = 8'h00;
    MEM[663] = 8'h00;
    MEM[664] = 8'h00;
    MEM[665] = 8'h00;
    MEM[666] = 8'h00;
    MEM[667] = 8'h00;
    MEM[668] = 8'h00;
    MEM[669] = 8'h00;
    MEM[670] = 8'h00;
    MEM[671] = 8'h00;
    MEM[672] = 8'h00;
    MEM[673] = 8'h00;
    MEM[674] = 8'h00;
    MEM[675] = 8'h00;
    MEM[676] = 8'h00;
    MEM[677] = 8'h00;
    MEM[678] = 8'h00;
    MEM[679] = 8'h00;
    MEM[680] = 8'h00;
    MEM[681] = 8'h00;
    MEM[682] = 8'h00;
    MEM[683] = 8'h00;
    MEM[684] = 8'h00;
    MEM[685] = 8'h00;
    MEM[686] = 8'h00;
    MEM[687] = 8'h00;
    MEM[688] = 8'h00;
    MEM[689] = 8'h00;
    MEM[690] = 8'h00;
    MEM[691] = 8'h00;
    MEM[692] = 8'h00;
    MEM[693] = 8'h00;
    MEM[694] = 8'h00;
    MEM[695] = 8'h00;
    MEM[696] = 8'h00;
    MEM[697] = 8'h00;
    MEM[698] = 8'h00;
    MEM[699] = 8'h00;
    MEM[700] = 8'h00;
    MEM[701] = 8'h00;
    MEM[702] = 8'h00;
    MEM[703] = 8'h00;
    MEM[704] = 8'h00;
    MEM[705] = 8'h00;
    MEM[706] = 8'h00;
    MEM[707] = 8'h00;
    MEM[708] = 8'h00;
    MEM[709] = 8'h00;
    MEM[710] = 8'h00;
    MEM[711] = 8'h00;
    MEM[712] = 8'h00;
    MEM[713] = 8'h00;
    MEM[714] = 8'h00;
    MEM[715] = 8'h00;
    MEM[716] = 8'h00;
    MEM[717] = 8'h00;
    MEM[718] = 8'h00;
    MEM[719] = 8'h00;
    MEM[720] = 8'h00;
    MEM[721] = 8'h00;
    MEM[722] = 8'h00;
    MEM[723] = 8'h00;
    MEM[724] = 8'h00;
    MEM[725] = 8'h00;
    MEM[726] = 8'h00;
    MEM[727] = 8'h00;
    MEM[728] = 8'h00;
    MEM[729] = 8'h00;
    MEM[730] = 8'h00;
    MEM[731] = 8'h00;
    MEM[732] = 8'h00;
    MEM[733] = 8'h00;
    MEM[734] = 8'h00;
    MEM[735] = 8'h00;
    MEM[736] = 8'h00;
    MEM[737] = 8'h00;
    MEM[738] = 8'h00;
    MEM[739] = 8'h00;
    MEM[740] = 8'h00;
    MEM[741] = 8'h00;
    MEM[742] = 8'h00;
    MEM[743] = 8'h00;
    MEM[744] = 8'h00;
    MEM[745] = 8'h00;
    MEM[746] = 8'h00;
    MEM[747] = 8'h00;
    MEM[748] = 8'h00;
    MEM[749] = 8'h00;
    MEM[750] = 8'h00;
    MEM[751] = 8'h00;
    MEM[752] = 8'h00;
    MEM[753] = 8'h00;
    MEM[754] = 8'h00;
    MEM[755] = 8'h00;
    MEM[756] = 8'h00;
    MEM[757] = 8'h00;
    MEM[758] = 8'h00;
    MEM[759] = 8'h00;
    MEM[760] = 8'h00;
    MEM[761] = 8'h00;
    MEM[762] = 8'h00;
    MEM[763] = 8'h00;
    MEM[764] = 8'h00;
    MEM[765] = 8'h00;
    MEM[766] = 8'h00;
    MEM[767] = 8'h00;
    MEM[768] = 8'h00;
    MEM[769] = 8'h00;
    MEM[770] = 8'h00;
    MEM[771] = 8'h00;
    MEM[772] = 8'h00;
    MEM[773] = 8'h00;
    MEM[774] = 8'h00;
    MEM[775] = 8'h00;
    MEM[776] = 8'h00;
    MEM[777] = 8'h00;
    MEM[778] = 8'h00;
    MEM[779] = 8'h00;
    MEM[780] = 8'h00;
    MEM[781] = 8'h00;
    MEM[782] = 8'h00;
    MEM[783] = 8'h00;
    MEM[784] = 8'h00;
    MEM[785] = 8'h00;
    MEM[786] = 8'h00;
    MEM[787] = 8'h00;
    MEM[788] = 8'h00;
    MEM[789] = 8'h00;
    MEM[790] = 8'h00;
    MEM[791] = 8'h00;
    MEM[792] = 8'h00;
    MEM[793] = 8'h00;
    MEM[794] = 8'h00;
    MEM[795] = 8'h00;
    MEM[796] = 8'h00;
    MEM[797] = 8'h00;
    MEM[798] = 8'h00;
    MEM[799] = 8'h00;
    MEM[800] = 8'h00;
    MEM[801] = 8'h00;
    MEM[802] = 8'h00;
    MEM[803] = 8'h00;
    MEM[804] = 8'h00;
    MEM[805] = 8'h00;
    MEM[806] = 8'h00;
    MEM[807] = 8'h00;
    MEM[808] = 8'h00;
    MEM[809] = 8'h00;
    MEM[810] = 8'h00;
    MEM[811] = 8'h00;
    MEM[812] = 8'h00;
    MEM[813] = 8'h00;
    MEM[814] = 8'h00;
    MEM[815] = 8'h00;
    MEM[816] = 8'h00;
    MEM[817] = 8'h00;
    MEM[818] = 8'h00;
    MEM[819] = 8'h00;
    MEM[820] = 8'h00;
    MEM[821] = 8'h00;
    MEM[822] = 8'h00;
    MEM[823] = 8'h00;
    MEM[824] = 8'h00;
    MEM[825] = 8'h00;
    MEM[826] = 8'h00;
    MEM[827] = 8'h00;
    MEM[828] = 8'h00;
    MEM[829] = 8'h00;
    MEM[830] = 8'h00;
    MEM[831] = 8'h00;
    MEM[832] = 8'h00;
    MEM[833] = 8'h00;
    MEM[834] = 8'h00;
    MEM[835] = 8'h00;
    MEM[836] = 8'h00;
    MEM[837] = 8'h00;
    MEM[838] = 8'h00;
    MEM[839] = 8'h00;
    MEM[840] = 8'h00;
    MEM[841] = 8'h00;
    MEM[842] = 8'h00;
    MEM[843] = 8'h00;
    MEM[844] = 8'h00;
    MEM[845] = 8'h00;
    MEM[846] = 8'h00;
    MEM[847] = 8'h00;
    MEM[848] = 8'h00;
    MEM[849] = 8'h00;
    MEM[850] = 8'h00;
    MEM[851] = 8'h00;
    MEM[852] = 8'h00;
    MEM[853] = 8'h00;
    MEM[854] = 8'h00;
    MEM[855] = 8'h00;
    MEM[856] = 8'h00;
    MEM[857] = 8'h00;
    MEM[858] = 8'h00;
    MEM[859] = 8'h00;
    MEM[860] = 8'h00;
    MEM[861] = 8'h00;
    MEM[862] = 8'h00;
    MEM[863] = 8'h00;
    MEM[864] = 8'h00;
    MEM[865] = 8'h00;
    MEM[866] = 8'h00;
    MEM[867] = 8'h00;
    MEM[868] = 8'h00;
    MEM[869] = 8'h00;
    MEM[870] = 8'h00;
    MEM[871] = 8'h00;
    MEM[872] = 8'h00;
    MEM[873] = 8'h00;
    MEM[874] = 8'h00;
    MEM[875] = 8'h00;
    MEM[876] = 8'h00;
    MEM[877] = 8'h00;
    MEM[878] = 8'h00;
    MEM[879] = 8'h00;
    MEM[880] = 8'h00;
    MEM[881] = 8'h00;
    MEM[882] = 8'h00;
    MEM[883] = 8'h00;
    MEM[884] = 8'h00;
    MEM[885] = 8'h00;
    MEM[886] = 8'h00;
    MEM[887] = 8'h00;
    MEM[888] = 8'h00;
    MEM[889] = 8'h00;
    MEM[890] = 8'h00;
    MEM[891] = 8'h00;
    MEM[892] = 8'h00;
    MEM[893] = 8'h00;
    MEM[894] = 8'h00;
    MEM[895] = 8'h00;
    MEM[896] = 8'h00;
    MEM[897] = 8'h00;
    MEM[898] = 8'h00;
    MEM[899] = 8'h00;
    MEM[900] = 8'h00;
    MEM[901] = 8'h00;
    MEM[902] = 8'h00;
    MEM[903] = 8'h00;
    MEM[904] = 8'h00;
    MEM[905] = 8'h00;
    MEM[906] = 8'h00;
    MEM[907] = 8'h00;
    MEM[908] = 8'h00;
    MEM[909] = 8'h00;
    MEM[910] = 8'h00;
    MEM[911] = 8'h00;
    MEM[912] = 8'h00;
    MEM[913] = 8'h00;
    MEM[914] = 8'h00;
    MEM[915] = 8'h00;
    MEM[916] = 8'h00;
    MEM[917] = 8'h00;
    MEM[918] = 8'h00;
    MEM[919] = 8'h00;
    MEM[920] = 8'h00;
    MEM[921] = 8'h00;
    MEM[922] = 8'h00;
    MEM[923] = 8'h00;
    MEM[924] = 8'h00;
    MEM[925] = 8'h00;
    MEM[926] = 8'h00;
    MEM[927] = 8'h00;
    MEM[928] = 8'h00;
    MEM[929] = 8'h00;
    MEM[930] = 8'h00;
    MEM[931] = 8'h00;
    MEM[932] = 8'h00;
    MEM[933] = 8'h00;
    MEM[934] = 8'h00;
    MEM[935] = 8'h00;
    MEM[936] = 8'h00;
    MEM[937] = 8'h00;
    MEM[938] = 8'h00;
    MEM[939] = 8'h00;
    MEM[940] = 8'h00;
    MEM[941] = 8'h00;
    MEM[942] = 8'h00;
    MEM[943] = 8'h00;
    MEM[944] = 8'h00;
    MEM[945] = 8'h00;
    MEM[946] = 8'h00;
    MEM[947] = 8'h00;
    MEM[948] = 8'h00;
    MEM[949] = 8'h00;
    MEM[950] = 8'h00;
    MEM[951] = 8'h00;
    MEM[952] = 8'h00;
    MEM[953] = 8'h00;
    MEM[954] = 8'h00;
    MEM[955] = 8'h00;
    MEM[956] = 8'h00;
    MEM[957] = 8'h00;
    MEM[958] = 8'h00;
    MEM[959] = 8'h00;
    MEM[960] = 8'h00;
    MEM[961] = 8'h00;
    MEM[962] = 8'h00;
    MEM[963] = 8'h00;
    MEM[964] = 8'h00;
    MEM[965] = 8'h00;
    MEM[966] = 8'h00;
    MEM[967] = 8'h00;
    MEM[968] = 8'h00;
    MEM[969] = 8'h00;
    MEM[970] = 8'h00;
    MEM[971] = 8'h00;
    MEM[972] = 8'h00;
    MEM[973] = 8'h00;
    MEM[974] = 8'h00;
    MEM[975] = 8'h00;
    MEM[976] = 8'h00;
    MEM[977] = 8'h00;
    MEM[978] = 8'h00;
    MEM[979] = 8'h00;
    MEM[980] = 8'h00;
    MEM[981] = 8'h00;
    MEM[982] = 8'h00;
    MEM[983] = 8'h00;
    MEM[984] = 8'h00;
    MEM[985] = 8'h00;
    MEM[986] = 8'h00;
    MEM[987] = 8'h00;
    MEM[988] = 8'h00;
    MEM[989] = 8'h00;
    MEM[990] = 8'h00;
    MEM[991] = 8'h00;
    MEM[992] = 8'h00;
    MEM[993] = 8'h00;
    MEM[994] = 8'h00;
    MEM[995] = 8'h00;
    MEM[996] = 8'h00;
    MEM[997] = 8'h00;
    MEM[998] = 8'h00;
    MEM[999] = 8'h00;
    MEM[1000] = 8'h00;
    MEM[1001] = 8'h00;
    MEM[1002] = 8'h00;
    MEM[1003] = 8'h00;
    MEM[1004] = 8'h00;
    MEM[1005] = 8'h00;
    MEM[1006] = 8'h00;
    MEM[1007] = 8'h00;
    MEM[1008] = 8'h00;
    MEM[1009] = 8'h00;
    MEM[1010] = 8'h00;
    MEM[1011] = 8'h00;
    MEM[1012] = 8'h00;
    MEM[1013] = 8'h00;
    MEM[1014] = 8'h00;
    MEM[1015] = 8'h00;
    MEM[1016] = 8'h00;
    MEM[1017] = 8'h00;
    MEM[1018] = 8'h00;
    MEM[1019] = 8'h00;
    MEM[1020] = 8'h00;
    MEM[1021] = 8'h00;
    MEM[1022] = 8'h00;
    MEM[1023] = 8'h00;
    MEM[1024] = 8'hfc;
    MEM[1025] = 8'hff;
    MEM[1026] = 8'hbd;
    MEM[1027] = 8'h23;
    MEM[1028] = 8'h00;
    MEM[1029] = 8'h00;
    MEM[1030] = 8'hbf;
    MEM[1031] = 8'haf;
    MEM[1032] = 8'ha5;
    MEM[1033] = 8'ha5;
    MEM[1034] = 8'h04;
    MEM[1035] = 8'h3c;
    MEM[1036] = 8'h5a;
    MEM[1037] = 8'h5a;
    MEM[1038] = 8'h84;
    MEM[1039] = 8'h34;
    MEM[1040] = 8'hac;
    MEM[1041] = 8'hac;
    MEM[1042] = 8'h05;
    MEM[1043] = 8'h20;
    MEM[1044] = 8'h0d;
    MEM[1045] = 8'h01;
    MEM[1046] = 8'h00;
    MEM[1047] = 8'h0c;
    MEM[1048] = 8'h02;
    MEM[1049] = 8'h00;
    MEM[1050] = 8'h40;
    MEM[1051] = 8'h1c;
    MEM[1052] = 8'had;
    MEM[1053] = 8'hde;
    MEM[1054] = 8'h10;
    MEM[1055] = 8'h20;
    MEM[1056] = 8'h0e;
    MEM[1057] = 8'h01;
    MEM[1058] = 8'h00;
    MEM[1059] = 8'h08;
    MEM[1060] = 8'h8e;
    MEM[1061] = 8'hd0;
    MEM[1062] = 8'h10;
    MEM[1063] = 8'h20;
    MEM[1064] = 8'h00;
    MEM[1065] = 8'h00;
    MEM[1066] = 8'hbf;
    MEM[1067] = 8'h8f;
    MEM[1068] = 8'h04;
    MEM[1069] = 8'h00;
    MEM[1070] = 8'hbd;
    MEM[1071] = 8'h23;
    MEM[1072] = 8'h08;
    MEM[1073] = 8'h00;
    MEM[1074] = 8'he0;
    MEM[1075] = 8'h03;
    MEM[1076] = 8'h00;
    MEM[1077] = 8'h43;
    MEM[1078] = 8'h04;
    MEM[1079] = 8'h00;
    MEM[1080] = 8'h04;
    MEM[1081] = 8'h48;
    MEM[1082] = 8'ha4;
    MEM[1083] = 8'h00;
    MEM[1084] = 8'ha5;
    MEM[1085] = 8'h55;
    MEM[1086] = 8'h0a;
    MEM[1087] = 8'h3c;
    MEM[1088] = 8'h00;
    MEM[1089] = 8'ha0;
    MEM[1090] = 8'h4a;
    MEM[1091] = 8'h35;
    MEM[1092] = 8'h01;
    MEM[1093] = 8'h00;
    MEM[1094] = 8'h48;
    MEM[1095] = 8'h11;
    MEM[1096] = 8'h27;
    MEM[1097] = 8'h01;
    MEM[1098] = 8'h00;
    MEM[1099] = 8'h08;
    MEM[1100] = 8'h01;
    MEM[1101] = 8'h00;
    MEM[1102] = 8'h49;
    MEM[1103] = 8'h11;
    MEM[1104] = 8'h27;
    MEM[1105] = 8'h01;
    MEM[1106] = 8'h00;
    MEM[1107] = 8'h08;
    MEM[1108] = 8'h02;
    MEM[1109] = 8'h43;
    MEM[1110] = 8'h04;
    MEM[1111] = 8'h00;
    MEM[1112] = 8'h06;
    MEM[1113] = 8'h48;
    MEM[1114] = 8'ha4;
    MEM[1115] = 8'h00;
    MEM[1116] = 8'h0a;
    MEM[1117] = 8'h00;
    MEM[1118] = 8'h0a;
    MEM[1119] = 8'h3c;
    MEM[1120] = 8'h55;
    MEM[1121] = 8'h5a;
    MEM[1122] = 8'h4a;
    MEM[1123] = 8'h35;
    MEM[1124] = 8'h01;
    MEM[1125] = 8'h00;
    MEM[1126] = 8'h48;
    MEM[1127] = 8'h11;
    MEM[1128] = 8'h27;
    MEM[1129] = 8'h01;
    MEM[1130] = 8'h00;
    MEM[1131] = 8'h08;
    MEM[1132] = 8'h01;
    MEM[1133] = 8'h00;
    MEM[1134] = 8'h49;
    MEM[1135] = 8'h11;
    MEM[1136] = 8'h27;
    MEM[1137] = 8'h01;
    MEM[1138] = 8'h00;
    MEM[1139] = 8'h08;
    MEM[1140] = 8'h03;
    MEM[1141] = 8'h43;
    MEM[1142] = 8'h04;
    MEM[1143] = 8'h00;
    MEM[1144] = 8'h07;
    MEM[1145] = 8'h48;
    MEM[1146] = 8'ha4;
    MEM[1147] = 8'h00;
    MEM[1148] = 8'hfa;
    MEM[1149] = 8'hff;
    MEM[1150] = 8'h0a;
    MEM[1151] = 8'h3c;
    MEM[1152] = 8'h55;
    MEM[1153] = 8'h5a;
    MEM[1154] = 8'h4a;
    MEM[1155] = 8'h35;
    MEM[1156] = 8'h01;
    MEM[1157] = 8'h00;
    MEM[1158] = 8'h48;
    MEM[1159] = 8'h11;
    MEM[1160] = 8'h27;
    MEM[1161] = 8'h01;
    MEM[1162] = 8'h00;
    MEM[1163] = 8'h08;
    MEM[1164] = 8'h01;
    MEM[1165] = 8'h00;
    MEM[1166] = 8'h49;
    MEM[1167] = 8'h11;
    MEM[1168] = 8'h27;
    MEM[1169] = 8'h01;
    MEM[1170] = 8'h00;
    MEM[1171] = 8'h08;
    MEM[1172] = 8'h01;
    MEM[1173] = 8'h00;
    MEM[1174] = 8'h02;
    MEM[1175] = 8'h24;
    MEM[1176] = 8'h08;
    MEM[1177] = 8'h00;
    MEM[1178] = 8'he0;
    MEM[1179] = 8'h03;
    MEM[1180] = 8'h21;
    MEM[1181] = 8'h10;
    MEM[1182] = 8'h00;
    MEM[1183] = 8'h00;
    MEM[1184] = 8'h08;
    MEM[1185] = 8'h00;
    MEM[1186] = 8'he0;
    MEM[1187] = 8'h03;

end
    
endmodule