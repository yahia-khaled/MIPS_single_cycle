module MIPS_single_cycle_tb();
    
endmodule