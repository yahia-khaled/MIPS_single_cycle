package MIPS_package;



endpackage